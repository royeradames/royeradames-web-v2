<svg xmlns="http://www.w3.org/2000/svg" width="4" height="100%" viewBox="0 0 4 100%" fill="none">
<rect x="0.5625" y="0.125" width="3" height="100%" fill="#ACB1C3"/>
</svg>
